library verilog;
use verilog.vl_types.all;
entity shiftrow_tb is
end shiftrow_tb;
