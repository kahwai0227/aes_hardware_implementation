library verilog;
use verilog.vl_types.all;
entity roundKeyGenerator_tb is
end roundKeyGenerator_tb;
