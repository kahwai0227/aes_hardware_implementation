library verilog;
use verilog.vl_types.all;
entity aes_testbench is
end aes_testbench;
