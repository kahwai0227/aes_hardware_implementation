library verilog;
use verilog.vl_types.all;
entity mixcolumn_tb is
end mixcolumn_tb;
