library verilog;
use verilog.vl_types.all;
entity aes_cudu_tb is
end aes_cudu_tb;
