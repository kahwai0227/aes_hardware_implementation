module mixColumns (
    input [7:0] state_matrix [0:3][0:3], // Input state matrix
    output reg [7:0] mixed_matrix [0:3][0:3] // Output mixed matrix
);

// Define the fixed matrix for MixColumns
reg [7:0] mix_matrix [0:3][0:3] = '{
    '{8'h02, 8'h03, 8'h01, 8'h01},
    '{8'h01, 8'h02, 8'h03, 8'h01},
    '{8'h01, 8'h01, 8'h02, 8'h03},
    '{8'h03, 8'h01, 8'h01, 8'h02}
};

// Perform MixColumns operation
always @* begin
    for (int col = 0; col < 4; col = col + 1) begin
        for (int row = 0; row < 4; row = row + 1) begin
            mixed_matrix[row][col] = 
                mix_column(state_matrix[0][col], state_matrix[1][col], state_matrix[2][col], state_matrix[3][col]);
        end
    end
end

// Function to perform the MixColumns operation for a single column
function [7:0] mix_column;
    input [7:0] a, b, c, d;
    begin
        case ({a, b, c, d})
            // Define multiplication in Galois Field (GF(2^8))
            8'h01: mix_column = a;
            8'h02: mix_column = a << 1;
            8'h03: mix_column = (a << 1) ^ a;
            default: mix_column = 8'h00; // For unused cases
        endcase
    end
endfunction

endmodule
