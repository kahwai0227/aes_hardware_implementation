library verilog;
use verilog.vl_types.all;
entity addRoundKey_tb is
end addRoundKey_tb;
