library verilog;
use verilog.vl_types.all;
entity aes_top_tb is
end aes_top_tb;
