library verilog;
use verilog.vl_types.all;
entity keyGenerator_tb is
end keyGenerator_tb;
