library verilog;
use verilog.vl_types.all;
entity rounds_tb is
end rounds_tb;
