library verilog;
use verilog.vl_types.all;
entity subbyte_tb is
end subbyte_tb;
