library verilog;
use verilog.vl_types.all;
entity aes_cu_tb is
end aes_cu_tb;
