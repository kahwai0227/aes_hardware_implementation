library verilog;
use verilog.vl_types.all;
entity mul_tb is
end mul_tb;
